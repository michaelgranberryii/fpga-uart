library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity fifo_ex_stat is
  generic(
     ADDR_WIDTH : integer := 2;
     DATA_WIDTH : integer := 8
  );
  port(
     clk, reset : in  std_logic;
     rd, wr     : in  std_logic;
     w_data     : in  std_logic_vector(DATA_WIDTH - 1 downto 0);
     empty      : out std_logic;
     full       : out std_logic;
     almost_empty, almost_full : out std_logic;
     word_count : out std_logic_vector(ADDR_WIDTH downto 0); 
     r_data     : out std_logic_vector(DATA_WIDTH - 1 downto 0)
  );
end fifo_ex_stat;

architecture Behavioral of fifo_ex_stat is
    signal full_tmp : std_logic;
    signal wr_en    : std_logic;
    signal w_addr   : std_logic_vector(ADDR_WIDTH - 1 downto 0);
    signal r_addr   : std_logic_vector(ADDR_WIDTH - 1 downto 0);

begin
-- write enabled only when FIFO is not full
  wr_en <= wr and (not full_tmp);
  full  <= full_tmp;
  
-- instantiate fifo control unit
  ctrl_unit : entity work.fifo_ctrl_ex_stat
     generic map(ADDR_WIDTH => ADDR_WIDTH)
     port map(
        clk    => clk,
        reset  => reset,
        rd     => rd,
        wr     => wr,
        empty  => empty,
        full   => full_tmp,
        almost_empty => almost_empty,
        almost_full => almost_full,
        word_count => word_count,
        w_addr => w_addr,
        r_addr => r_addr);
        
-- instantiate register file
  reg_file_unit : entity work.reg_file
     generic map(
        DATA_WIDTH => DATA_WIDTH,
        ADDR_WIDTH => ADDR_WIDTH)
     port map(
        clk    => clk,
        w_addr => w_addr,
        r_addr => r_addr,
        w_data => w_data,
        r_data => r_data,
        wr_en  => wr_en);

end Behavioral;
